library verilog;
use verilog.vl_types.all;
entity conv_kernel_tb is
end conv_kernel_tb;
